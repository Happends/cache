module test;

    cache cache();
    intial begin
        #1;
        $finsish;
endmodule